--/*
--  *******************************************************
--  Computer Architecture Course, Laboratory Sources 
--  Amirkabir University of Technology (Tehran Polytechnic)
--  Department of Computer Engineering (CE-AUT)
--  https://ce[dot]aut[dot]ac[dot]ir
--  Designed by Ali Mohammadpour(@alimpk)
--  *******************************************************
--  All Rights reserved (C) 2019-2020
--  *******************************************************
--  Student ID  : 
--  Student Name: 
--  Student Mail: 
--  *******************************************************
--  Additional Comments:
--
--*/

-----------------------------------------------------------
---  Module Name: Ripple Counter 
---  Description: 4 Bit Ripple Counter
-----------------------------------------------------------
entity ripple_counter is

	port (
		clk     : in  std_logic;
		rst     : in  std_logic;
		count : out std_logic_vector(3 downto 0)
	);
end ripple_counter;

architecture comprator_arc of ripple_counter is
begin
signal wire : std_logic_vector(9 downto 0)
First_TFF : 



end comprator_arc;
